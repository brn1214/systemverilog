class cfg;
    // Integer fields with default values
    int latency = 1; // 'latency' field with a default value of 1.
    int amount = 10; // 'amount' field with a default value of 10.

endclass
